package moore_pack is                			-- Декларация пакета
	type state_s is (a1,a2,a3,a4,a5,a6);		-- Алфавит состояний
end package moore_pack;
